`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/11/12 15:58:19
// Design Name: 
// Module Name: alu_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu_tb;
reg [31:0]a;
reg [31:0]b;
reg [3:0]aluc;
wire [31:0]r;
wire zero;
wire carry;
wire negative;
wire overflow;
alu uut (.a(a),
.b(b),
.aluc(aluc),
.r(r),
.zero(zero),
.carry(carry),
.negative(negative),
.overflow(overflow));

initial
begin
aluc=4'b0000;
    a=0;
    b=0;
    #10
    a=0;
    b=1;
    #10
    a={32{1'b1}};
    b=1;
    #10
    a={32{1'b1}};
    b={32{1'b1}};
     #10                 
    a={1'b0,{31{1'b1}}};
    b={1'b0,{31{1'b1}}};
    #50
    
    aluc=4'b0010;
    a=0;
    b=0;
    #10
    a=0;
    b=1;
    #10
    a={32{1'b1}};
    b=1;
    #10
    a={32{1'b1}};
    b={32{1'b1}};
    #10
    a={1'b0,{31{1'b1}}};
    b={1'b0,{31{1'b1}}};
    #50
    
    aluc=4'b0001;
    a=0;
    b=0;
    #10
    a=0;
    b=1;
    #10
    a={32{1'b1}};
    b=1;
    #10
    a={32{1'b1}};
    b={32{1'b1}};
     #10                 
    a={1'b0,{31{1'b1}}};
    b={1'b0,{31{1'b1}}};
    #50
    
      aluc=4'b0011;
      a=0;
      b=0;
      #10
      a=0;
      b=1;
      #10
      a={32{1'b1}};
      b=1;
      #10
      a={32{1'b1}};
      b={32{1'b1}};
      #10
      a={1'b0,{31{1'b1}}};
      b={1'b0,{31{1'b1}}};
     #10
     a={1'b0,{31{1'b1}}};
     b={1'b1,{31{1'b1}}};
    
     aluc=4'b0100;
     a={{8{1'b1}},{8{1'b0}},{8{1'b0}},{8{1'b1}}};
     b={{8{1'b1}},{8{1'b1}},{8{1'b0}},{8{1'b0}}};
     #10
     aluc=4'b0101;
     a={{8{1'b1}},{8{1'b0}},{8{1'b0}},{8{1'b1}}};
     b={{8{1'b1}},{8{1'b1}},{8{1'b0}},{8{1'b0}}};
     #10
     aluc=4'b0110;
     a={{8{1'b1}},{8{1'b0}},{8{1'b0}},{8{1'b1}}};
     b={{8{1'b1}},{8{1'b1}},{8{1'b0}},{8{1'b0}}};
     #10
     aluc=4'b0111;
     a={{8{1'b1}},{8{1'b0}},{8{1'b0}},{8{1'b1}}};
     b={{8{1'b1}},{8{1'b1}},{8{1'b0}},{8{1'b0}}};
     
    aluc =4'b1000;
     b={{16{1'b0}},{16{1'b1}}};
     #10
     aluc =4'b1001;
     b={{16{1'b1}},{16{1'b0}}};
     
     aluc = 4'b1011;
     a={1'b1,{31{1'b0}}};
     b={1'b0,{31{1'b1}}};
     #10
     aluc = 4'b1010;
     
   aluc=4'b1100;
    b={1'b0,{31{1'b1}}};
    a=32'd32;
    #10
    b={1'b1,{31{1'b0}}};
    a=32'd32;
    #10
    b=32'b101010;
    a=32'd3;
    aluc=4'b1101;
    b={1'b0,{31{1'b1}}};
    a=32'd32;
    #10
    b={1'b1,{31{1'b0}}};
    a=32'd32;
    #10
    b=32'b101010;
    a=32'd3;
    
    aluc=4'b1111;
     b={16'b0,{16{1'b1}}};
     a=32'd16;
     #10
     b={16'b1,{16{1'b0}}};
     a=32'd16;

end
endmodule
